module TRNG (
    input wire clk,
    input wire rst_n,

    input wire trng_request,
    output wire [31:0] random_number,
    output wire ready
);

    // TRNG implementation goes here

endmodule
