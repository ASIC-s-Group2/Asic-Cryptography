module CC20TopLevel(
    input wire clk,
    input wire reset,
    input wire [255:0] key,
    input wire [127:0] plaintext,
)
endmodule
